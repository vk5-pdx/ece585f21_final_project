/****************************************************************
 * queue_tb.sv - testbench for queue
 *
 * Author        : Viraj Khatri (vk5@pdx.edu)
 * Last Modified : 16th November, 2021
 *
 * Description   :
 * -----------
 * testbench for queue
 ****************************************************************/

module queue_tb;

logic clk, rst_n;

endmodule : queue_tb
